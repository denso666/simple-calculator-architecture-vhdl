library ieee;
use ieee.std_logic_1164.all;

entity test_bench is end entity;

architecture behavior of test_bench is begin

end architecture;